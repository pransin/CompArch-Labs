module shifter(in, pc, out);
input [26:0]in;
input [4:0]pc
output
endmodule