module pc(out, in);
input [4:0] in;
output reg[4:0] out;

endmodule