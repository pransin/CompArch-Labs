module test_bench(clk, rst);
  input  clk;
  input  rst;
  wire   [31:0] wire_39069600;
  wire   [31:0] wire_39795024;
  wire   [31:0] wire_39795168;
  wire   wire_39795168_stb;
  file_reader_a file_reader_a_39796104(
    .clk(clk),
    .rst(rst),
    .AbyB(wire_39069600),
    .DONE(wire_39069600_stb),
  file_reader_b file_reader_b_39759816(
    .clk(clk),
    .rst(rst),
    .AbyB(wire_39795024),
    .DONE(wire_39795024_stb),
  file_writer file_writer_39028208(
    .clk(clk),
    .rst(rst),
    .input_a(wire_39795168),
  divider divider_39759952(
    .clk(clk),
    .rst(rst),
    .input_a(wire_39069600),
    .input_a_stb(wire_39069600_stb),
    .input_a_ack(wire_39069600_ack),
    .input_b(wire_39795024),
    .input_b_stb(wire_39795024_stb),
    .input_b_ack(wire_39795024_ack),
    .output_z(wire_39795168),
    .output_z_stb(wire_39795168_stb),
    .output_z_ack(wire_39795168_ack));
endmodule